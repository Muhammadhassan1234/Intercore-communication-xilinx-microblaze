// -------------------------------------------------------------------------------------------------
// Designer:
// Description: 
// -------------------------------------------------------------------------------------------------

// -------------------------------------------------------------------------------------------------
// Module definition
// -------------------------------------------------------------------------------------------------
module module_name #(
  parameter RESET_ACTIVE_VALUE
) (
  input logic clk,
  input logic rst,
);

  // ---------------------------------------------------------------------------------------------
  // Declarations of the module_name
  // ---------------------------------------------------------------------------------------------

  // ---------------------------------------------------------------------------------------------
  // Implementation of the module_name
  // ---------------------------------------------------------------------------------------------

endmodule : module_name